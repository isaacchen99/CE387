    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.dropbox.attrs    

�=XwA��     L���ö�