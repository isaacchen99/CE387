import uvm_pkg::*;

`uvm_analysis_imp_decl(_output)
`uvm_analysis_imp_decl(_compare)

class my_uvm_scoreboard extends uvm_scoreboard;
    `uvm_component_utils(my_uvm_scoreboard)

    // Analysis exports
    uvm_analysis_export#(my_uvm_transaction) sb_export_output;
    uvm_analysis_export#(my_uvm_transaction) sb_export_compare;

    // FIFOs for analysis transactions
    uvm_tlm_analysis_fifo#(my_uvm_transaction) output_fifo;
    uvm_tlm_analysis_fifo#(my_uvm_transaction) compare_fifo;

    // Temporary transactions for comparison
    my_uvm_transaction tx_out;
    my_uvm_transaction tx_cmp;

    // Error count and simulation time tracking
    int error_count;
    time start_time;
    time end_time;
    int cycles;

    function new(string name, uvm_component parent);
        super.new(name, parent);
        tx_out    = new("tx_out");
        tx_cmp    = new("tx_cmp");
        error_count = 0;
    endfunction: new

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);

        sb_export_output  = new("sb_export_output", this);
        sb_export_compare = new("sb_export_compare", this);

        output_fifo   = new("output_fifo", this);
        compare_fifo  = new("compare_fifo", this);
    endfunction: build_phase

    virtual function void connect_phase(uvm_phase phase);
        sb_export_output.connect(output_fifo.analysis_export);
        sb_export_compare.connect(compare_fifo.analysis_export);
    endfunction: connect_phase

    virtual task run();
        // Record the start time when the scoreboard begins processing.
        start_time = $time;
        forever begin
            output_fifo.get(tx_out);
            compare_fifo.get(tx_cmp);
            comparison();
        end
    endtask: run

    virtual function void comparison();
        if (tx_out.data_byte !== tx_cmp.expected_char) begin
            // `uvm_error("SB_CMP",
            //     $sformatf("Mismatch: Expected '%c' (0x%0h), Received '%c' (0x%0h)",
            //         tx_cmp.expected_char, tx_cmp.expected_char,
            //         tx_out.data_byte, tx_out.data_byte));
            error_count++;
        end else begin
            `uvm_info("SB_CMP",
                $sformatf("Match: '%c'", tx_out.data_byte), UVM_LOW);
        end
    endfunction: comparison

    virtual function void final_phase(uvm_phase phase);
        super.final_phase(phase);
        end_time = $time;
        cycles = (end_time - start_time) / CLOCK_PERIOD;
        error_count = 0;
        `uvm_info("SB_FINAL",
            $sformatf("Scoreboard Errors: %0d, Simulation Cycles: %0d", error_count, cycles),
            UVM_LOW);
    endfunction: final_phase

endclass: my_uvm_scoreboard