package my_uvm_package;

import uvm_pkg::*;

// UVM files
`include "uvm_macros.svh"
`include "my_uvm_transaction.sv"
`include "my_uvm_globals.sv"
`include "my_uvm_sequence.sv"
`include "my_uvm_monitor.sv"
`include "my_uvm_driver.sv"
`include "my_uvm_agent.sv"
`include "my_uvm_scoreboard.sv"
`include "my_uvm_config.sv"
`include "my_uvm_env.sv"
`include "my_uvm_test.sv"

endpackage
