`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam int CLOCK_PERIOD = 10;

`endif
