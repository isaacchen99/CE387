module udp_parser_top (
  input  logic         clk,
  input  logic         reset,
  // Testbench input interface: stream a UDP packet (with SOF/EOF markers)
  input  logic [7:0]   tb_in_data,
  input  logic         tb_in_valid,
  input  logic         tb_in_sof,
  input  logic         tb_in_eof,
  output logic         tb_in_ready,
  // Testbench output interface: read the decoded UDP payload
  output logic [7:0]   tb_out_data,
  output logic         tb_out_valid,
  output logic         tb_out_sof,
  output logic         tb_out_eof,
  input  logic         tb_out_ready
);

  //-------------------------------------------------------------------------
  // Wires connecting the input ctrl_fifo to the UDP parser
  //-------------------------------------------------------------------------
  wire [7:0] in_fifo_rdata;
  wire       in_fifo_rvalid;
  wire       in_fifo_rsof;
  wire       in_fifo_reof;
  // When the input FIFO is empty, r_valid is low.
  wire       in_fifo_empty = ~in_fifo_rvalid;
  
  // This signal is generated by the UDP parser to tell the input FIFO when it’s ready
  wire       parser_in_ready;
  
  //-------------------------------------------------------------------------
  // Instantiate the input FIFO controller.
  // This FIFO accepts the framed UDP packet from the testbench.
  //-------------------------------------------------------------------------
  ctrl_fifo in_ctrl_fifo_inst (
    .clk    (clk),
    .reset  (reset),
    // Write side driven by testbench
    .wdata  (tb_in_data),
    .w_valid(tb_in_valid),
    .w_sof  (tb_in_sof),
    .w_eof  (tb_in_eof),
    .w_ready(tb_in_ready),
    // Read side drives the UDP parser
    .rdata  (in_fifo_rdata),
    .r_valid(in_fifo_rvalid),
    .r_sof  (in_fifo_rsof),
    .r_eof  (in_fifo_reof),
    .r_ready(parser_in_ready)
  );
  
  //-------------------------------------------------------------------------
  // Wires connecting the UDP parser to the output FIFO controller.
  //-------------------------------------------------------------------------
  wire [7:0] parser_out_data;
  wire       parser_out_valid;
  wire       parser_out_sof;
  wire       parser_out_eof;
  
  // The UDP parser’s output ready is driven by the output FIFO’s ability
  // to accept new data. (We derive out_fifo_full from the output FIFO's write-ready.)
  wire       out_fifo_wready;
  wire       out_fifo_full = ~out_fifo_wready;
  // The UDP parser's out_ready signal is the same as the output FIFO's write ready.
  wire       parser_out_ready;
  assign parser_out_ready = out_fifo_wready;
  
  // For debugging/error reporting from the UDP parser.
  wire       parser_error_flag;
  
  //-------------------------------------------------------------------------
  // Instantiate the UDP parser.
  // The UDP parser reads from the input FIFO and streams out the decoded UDP payload.
  //-------------------------------------------------------------------------
  udp_parser udp_parser_inst (
    .clk            (clk),
    .rst_n          (~reset),
    // Input side (from in_ctrl_fifo)
    .in_data        (in_fifo_rdata),
    .in_valid       (in_fifo_rvalid),
    .in_sof         (in_fifo_rsof),
    .in_eof         (in_fifo_reof),
    .in_fifo_empty  (in_fifo_empty),
    .in_ready       (parser_in_ready),
    // Output side (to out_ctrl_fifo)
    .out_data       (parser_out_data),
    .out_valid      (parser_out_valid),
    .out_sof        (parser_out_sof),
    .out_eof        (parser_out_eof),
    .out_ready      (parser_out_ready),
    .out_fifo_full  (out_fifo_full),
    .error_flag     (parser_error_flag)
  );
  
  //-------------------------------------------------------------------------
  // Instantiate the output FIFO controller.
  // This FIFO collects the decoded UDP payload from the UDP parser and
  // presents it (with new SOF/EOF markers) to the testbench.
  //-------------------------------------------------------------------------
  ctrl_fifo out_ctrl_fifo_inst (
    .clk    (clk),
    .reset  (reset),
    // Write side driven by UDP parser output
    .wdata  (parser_out_data),
    .w_valid(parser_out_valid),
    .w_sof  (parser_out_sof),
    .w_eof  (parser_out_eof),
    .w_ready(out_fifo_wready),
    // Read side driven by testbench
    .rdata  (tb_out_data),
    .r_valid(tb_out_valid),
    .r_sof  (tb_out_sof),
    .r_eof  (tb_out_eof),
    .r_ready(tb_out_ready)
  );
  
endmodule